------------------------------------------------------------------------------
-- This file is part of 'SLAC EVR Gen2'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'SLAC EVR Gen2', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package Version is

   constant FPGA_VERSION_C : std_logic_vector(31 downto 0) := x"CED20020";  -- MAKE_VERSION

   constant BUILD_STAMP_C : string := "LegacyEvrCardG2: Vivado v2015.4 (x86_64) Built Fri Apr 15 16:10:24 PDT 2016 by ruckman";

end Version;

-------------------------------------------------------------------------------
-- Revision History:
--
-- 07/24/2015 (CED20000): Initial Build
-- 07/30/2015 (CED20001): Inverted the output to match Legacy EVR output
-- 08/06/2015 (CED20002): In getPcieHdr(), reordered FirstDwBe & LastDwBe
-- 08/17/2015 (CED20003): Fixed the 16-bit accesses in the EvrV1Reg.vhd
-- 08/17/2015 (CED20004): Fixed the intFlag(3) importing bug
-- 08/18/2015 (CED20005): In EvrV1TimeStampFIFO.vhd, change FWFT_EN_G from "false" to "true"
-- 09/23/2015 (CED20006): Removed 4 shift registers in EvrV1EventReceiver for rxData & rxDataK
--                        Registering the trigger outputs and set the SLEW = FAST
-- 09/24/2015 (CED20007): Added 2 cycles address setup delay for BRAM's AXI-Lite read transactions
-- 09/25/2015 (CED20008): Removed the dbRdAddr Synchronizer 
--                        Note: In EvrCardG2Trig.vhd: ODDR = "OPPOSITE_EDGE"
-- 10/19/2015 (CED20009): In EvrCardG2Trig.vhd: ODDR = "SAME_EDGE" and with clock MUX
-- 10/19/2015 (CED2000A): In EvrCardG2Trig.vhd: ODDR = "SAME_EDGE" and bypass clock MUX
-- 10/26/2015 (CED2000B): 
--    Revision Control:    Branching from CED2000A
--    In EVR core,         If no heartbeat event is received the counter times out (approx. 1.6 s)
--                         and a heartbeat flag is set.
--
-- 10/27/2015 (CED2000C): 
--    Revision Control:    Branching from CED2000B
--    In EVR core,         Synchronizing all status bits used to generate an interrupt on the axiClk
--                         clock domain and no longer a mix of axiClk/evrClk domain.
--
-- 10/28/2015 (CED2000D): 
--    Revision Control:    Branching from CED2000C
--    In EVR core,         Changed the Output Trigger Crossbar from registered to combinatory 
--                         to phase match with the MRF (removes 8.4 ns delay)
--    In MGT core,         If linkDown then, forward rxData = 0x0 and rxDataK = 0x0 to EVR core
--    In EvrCardG2Trig,    Bypass the trig MUX
--
-- 03/15/2016 (CED2000E): 
--    Revision Control:    Branching from CED2000D
--    In Top Level ,       Rebuilding the baseline 
--
-- 03/15/2016 (CED2000F): 
--    Revision Control:    Branching from CED2000E
--    In Top Level ,       Changed BPI from ASYNC to SYNC mode (TYPE2) and config clock from 9 MHz to 50 MHz 
--
-- 03/25/2016 (CED20010): 
--    Revision Control:    Branching from CED2000F
--    In Top Level ,       Disabled the ability for AxiVersion to cause a reboot of FPGA via PCIe register transaction
--
-- 04/04/2016 (CED20011): 
--    Revision Control:    Branching from CED20010
--    In PCI core,         Upgrade the Xilinx PCIe IP core from version 3.1 to version 3.2
--
-- 04/04/2016 (CED20012): 
--    Revision Control:    Branching from CED20011
--    In PCI core,         Debouncing the PCIe's reset for 1.5 us
--
-- 04/04/2016 (CED20013): 
--    Revision Control:    Branching from CED20012
--    In PCI core,         Debouncing the PCIe's reset for 10 ms
--
-- 04/05/2016 (CED20014): 
--    Revision Control:    Branching from CED20013
--    In PCI core,         Removed the debouncer (it didn't help or make worse the enumeration issue)
--    In PCI core,         Change the IP core to 
--                            1) c_disable_tx_aspm_l0s = TRUE
--                            2) c_ep_l0s_accpt_lat = 0
--                            3) ep_l0s_accpt_lat = 111
--                            4) Acceptable_L0s_Latency = Maximum_of_64_ns
--
-- 04/05/2016 (CED20015): 
--    Revision Control:    Branching from CED20014
--    In top level,        Terminating the unused PGP GT-CLK port
--
-- 04/06/2016 (CED20016): 
--    Revision Control:    Branching from CED20011
--    In top level,        Terminating the unused PGP GT-CLK port
--
-- 04/07/2016 (CED20017): 
--    Revision Control:    Branching from CED20010
--    In EVR core,         Added the following registers (based on Figure 1 of EVR-MRM-006.doc on page 7)
--                            0x05C    SecSR          UINT32   Seconds Shift Register
--                            0x060    SecCounter     UINT32   Timestamp Seconds Counter
--                            0x064    EventCounter   UINT32   Timestamp Event Counter
--                            0x068    SecLatch       UINT32   Timestamp Seconds Counter Latch
--                            0x06C    EvCntLatch     UINT32   Timestamp Event Counter Latch
--    In EVR core,         r.controlReg(9) is auto-clear in firmware
--    In EVR core,         r.controlReg(9) is used to latch the values for SecLatch & EvCntLatch
--    In Top Level,        Enable the ability for AxiVersion to cause a reboot of FPGA via PCIe register transaction
--                         Note: This ability is required for reloading the FPGA firmware without a cold reboot.
--
-- 04/07/2016 (CED20018): 
--    Revision Control:    Branching from CED20017
--    In EVR core,         Changed config.latchTs from r.controlReg(9) to r.controlReg(10)
--
-- 04/08/2016 (CED20019): 
--    Revision Control:    Branching from CED20018
--    In EVR core,         Added EvrCardG2LclsV1LedRgb.vhd
--
-- 04/08/2016 (CED2001A): 
--    Revision Control:    Branching from CED20019
--    In Common core,      Increase stable link status wait time from 0xFF to 0xFFFF (EvrGtp7.vhd's cnt)
--                         Changed gtRxResetDone from SYNC reset to ASYNC reset for stable link status
--                         Using the PCIe clock as stable reference, which prevents an oscillating state of 
--                         locked to not locked when establishing a new link.
--
-- 04/08/2016 (CED2001B): 
--    Revision Control:    Branching from CED2001A
--    In EVR core,         In EvrCardG2LclsV1LedRgb.vhd, registering the opCodeDet before going into a ASYNC reset port
--    In PCI core,         Upgrade the Xilinx PCIe IP core from version 3.1 to version 3.2
--    In PCI core,         Change the following PCIe PHY properties:
--                            1) In Capabilities[48]: 
--                               Changed from "64bit-" to "64bit+"
--                            2) In Capabilities[60].DevCap: 
--                               Changed from "Latency L0s unlimited, L1 unlimited" to "Latency L0s <64ns, L1 <1us"
--                            3) In Capabilities[60].DevCap2: 
--                               Changed from "Completion Timeout: Range B" to "Completion Timeout: Range A"
--
-- 04/12/2016 (CED2001C): 
--    Revision Control:    Branching from CED2001B
--    In EVR core,         Auto-reset the irqClear bus to 0x0 after register write
--
-- 04/12/2016 (CED2001D): 
--    Revision Control:    Branching from CED2001C
--    In EVR core,         In software (based on EVR-MRM-006.doc), the order of event FIFO readouts is:
--                            1) 0x78 event code (first read)
--                            2) 0x70 second register
--                            3) 0x74 timestamp register (last read)
--                         which is why the read FIFO strobe that's automatically generated from a read register 
--                         transaction was moved from ReadAddress@0x78 to ReadAddress@0x74
--
-- 04/12/2016 (CED2001E): 
--    Revision Control:    Branching from CED2001D
--    In Top Level ,       Disabled the ability for AxiVersion to cause a reboot of FPGA via PCIe register transaction
--    In EVR core,         Block all read transactions for 512 ns after set to r.controlReg(10) = 0x1 to 
--                         compensate for the latency of latching the time stamp bus
--                         Note: 512 ns is not an optimized value
--
-- 04/13/2016 (CED2001F): 
--    Revision Control:    Branching from CED2001E
--    In EVR core,         Optimized the block of all read transactions after r.controlReg(10) = 0x1 to 128 ns
--
-- 04/15/2016 (CED20020): 
--    Revision Control:    Branching from CED2001F
--    In TOP core,         Adding YAML support for firmware register definition (work in progress)
--
-------------------------------------------------------------------------------
